`timescale 1ns/10ps


module fifo_async_circular_tb ();



endmodule