`timescale 1ns/10ps


module fifo_tb ();



endmodule
